module and_gate(input1, input2, output_data);
    input input1, input2;
    output output_data;

    assign output_data = input1 & input2;
endmodule
